library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity DispCntrl is
	port(
	
	
	);
end DispCntrl;


architecture FSM of DispCntrl is
	

end FSM;